module diff_out (
		input  wire [0:0] din,       //       din.export
		output wire [0:0] pad_out,   //   pad_out.export
		output wire [0:0] pad_out_b  // pad_out_b.export
	);
endmodule

