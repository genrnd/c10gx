module sfl (
		input  wire  noe_in  // noe_in.noe
	);
endmodule

