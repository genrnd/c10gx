module diff_in (
		output wire [0:0] dout,     //     dout.export
		input  wire [0:0] pad_in,   //   pad_in.export
		input  wire [0:0] pad_in_b  // pad_in_b.export
	);
endmodule

